// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module objects_rom
   (
	 input wire clk,
    input wire [7:0] addr,
    output reg [31:0] data
   );

	/* Signal declaration */
   reg [7:0] addr_reg; 

   always @(posedge clk) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)
			
         //LETALO voznik
			8'h00: data = 32'b00000000000000000000000000000000; // 
			8'h01: data = 32'b00000000000000000000000000000000; // 
         8'h02: data = 32'b00000000000000011000000000000000; // 
			8'h03: data = 32'b00000000000000111100000000000000; // 
			8'h04: data = 32'b00000000000001111110000000000000; // 
			8'h05: data = 32'b00000000000001111110000000000000; // 
			8'h06: data = 32'b00000000000001111110000000000000; // 
			8'h07: data = 32'b00000000000001111110000000000000; // 
			8'h08: data = 32'b00000000000001111110000000000000; // 
			8'h09: data = 32'b00000000000001111110000000000000; // 
			8'h0a: data = 32'b00000000000011111111000000000000; // 
			8'h0b: data = 32'b00000000000011111111000000000000; //
			8'h0c: data = 32'b00000000000011111111000000000000; //
			8'h0d: data = 32'b00000000000001111110000000000000; // 
			8'h0e: data = 32'b00000001100100111100100110000000; // 
			8'h0f: data = 32'b00000011101111111111110111000000; // 
			8'h10: data = 32'b00001111111110111101111111110000; // 
			8'h11: data = 32'b00001111011110111101111011110000; // 
			8'h12: data = 32'b00111111000110111101100011111100; // 
			8'h13: data = 32'b01111111110110111101101111111110; // 
			8'h14: data = 32'b01111111011110111101111011111110; // 
			8'h15: data = 32'b11111111001110111101110011111111; // 
			8'h16: data = 32'b11111000000010111101000000011111; // 
			8'h17: data = 32'b11000000000111111111100000000011; // 
			8'h18: data = 32'b00000000001111111111110000000000; // 
			8'h19: data = 32'b00000000000111111111100000000000; // 
			8'h1a: data = 32'b00000000000000111100000000000000; // 
			8'h1b: data = 32'b00000000000011111111000000000000; // 
			8'h1c: data = 32'b00000000000111111111100000000000; // 
			8'h1d: data = 32'b00000000000110011001100000000000; // 
			8'h1e: data = 32'b00000000000000000000000000000000; // 
			8'h1f: data = 32'b00000000000000000000000000000000; // 


			// LETALO nasprotnik
         8'h20: data = 32'b00000000000011100111000000000000;
			8'h21: data = 32'b00000000000011111111000000000000;
			8'h22: data = 32'b00000000011111111111111000000000;
			8'h23: data = 32'b00011111111111111111111111111000;
			8'h24: data = 32'b01111111111111111111111111111110;
			8'h25: data = 32'b01111111111111111111111111111110;
			8'h26: data = 32'b01111111111111111111111111111110;
			8'h27: data = 32'b01111111111111100111111111111110;
			8'h28: data = 32'b01111111111111100111111111111110;
			8'h29: data = 32'b00111110111111100111111101111110;
			8'h2a: data = 32'b00011110011111100111111001111000;
			8'h2b: data = 32'b00000000011111100111111000000000;
			8'h2c: data = 32'b00000000001111100111110000000000;
			8'h2d: data = 32'b00000000001111111111110000000000;
			8'h2e: data = 32'b00000000001111111111110000000000;
			8'h2f: data = 32'b00000000001111111111110000000000;
			8'h30: data = 32'b00000000000011111111000000000000;
			8'h31: data = 32'b00000000000011111111000000000000;
			8'h32: data = 32'b00000000000011111111000000000000;
			8'h33: data = 32'b00000000000111111111100000000000;
			8'h34: data = 32'b00000000000111111111100000000000;
			8'h35: data = 32'b00000000000111111111100000000000;
			8'h36: data = 32'b00000000000110111101100000000000;
			8'h37: data = 32'b00000000000111111111100000000000;
			8'h38: data = 32'b00000000000111111111100000000000;
			8'h39: data = 32'b00000000000011111111000000000000;
			8'h3a: data = 32'b00000000000011111111000000000000;
			8'h3b: data = 32'b00000000000001111110000000000000;
			8'h3c: data = 32'b00000000000001111110000000000000;
			8'h3d: data = 32'b00000000000000111100000000000000;
			8'h3e: data = 32'b00000000000000111100000000000000;
			8'h3f: data = 32'b00000000000000011000000000000000;



			// STREL
			8'h40: data = 32'b00000000000000011000000000000000; // 
			8'h41: data = 32'b00000000000000111100000000000000; // 
			8'h42: data = 32'b00000000000000111100000000000000; // 
			8'h43: data = 32'b00000000000000111100000000000000; // 
			8'h44: data = 32'b00000000000000111100000000000000; // 
			8'h45: data = 32'b00000000000000111100000000000000; // 
			8'h46: data = 32'b00000000000000011000000000000000; // 

			default: data = 0;
   endcase  
   	       
endmodule      
	       
	       
	       
	       
	       
	       
	       